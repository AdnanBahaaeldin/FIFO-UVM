package FIFO_Shared_pkg;

//Define the FIFO_WIDTH and FIFO_DEPTH parameters
parameter FIFO_WIDTH = 16;
parameter FIFO_DEPTH = 8;

//Define Error and correct count variables
integer error_count, correct_count;

endpackage




